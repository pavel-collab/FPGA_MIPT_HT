/*
В книге А. Л. Ларина "Основы цифровой электроники" писаны 2 варианта реализации SR защелок --
на логическом "И" и на логическом "ИЛИ". Так как временные диаграммы приведены для защелки на 
логическом "ИЛИ", а в составе D защелок используется реализация на логическом "И",
в текущей дериктории представлены две реализации SR защелки
SR_OR_Latch.v -- на логическом "ИЛИ"
SR_Latch.v -- на логическом "И"
*/
// S, R -- входные шины, C -- шина состояния
module SR_Latch(
    input wire S, // Set
    input wire R, // Reset
    input wire C, // Condition
    output wire Q,
    output wire nQ
);
    assign Q = (~(R & nQ)&C);
    assign nQ = (~(S & Q)&C);

endmodule